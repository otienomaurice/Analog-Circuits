This is a ac sweep analysis of the circuit given
R1 1 2 10K;
R2 2 0 10K;
R3 2 3 10K;
R4 3 0 10K;
R5 3 4 10K;
C  4 0 0.01uF;
Vsig 1 0 DC 5v AC 1;
.AC DEC 20 10 100k;
.Probe;
.end;
