*Amplifier simulation

* Example of Amplifier Subcircuit instantiation and test
* Filename: Amplifier_test.cir,  Subcircuit called: Amplifier,  Subcircuit Definition file: Amplifier.sub

* Input Voltage source and resistance
Vsig 1 0 DC 0V AC 1v
R1 1 2 10K

* Load Resistance
Rload 3 0 1K

* Subcircuit instantiation.  All subcircuits start with leading character X and then unique identifier.
* Note:  The PINS must be in the correct order to match that of the subcircuit.
* In this case 2 = VIN  3 = VOUT and 0 = VGND  which matches order in sub file .subckt command.
Xamp 2 3 0 Amplifier

* Include card tells Spice to pull named file into this deck
.include Amplifier.sub

*Usual Spice Simulation Commands
.Ac DEC 20 1 1000000
.probe
.end

